library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.finish;
use work.all;

entity registro_32x32_tb is
end registro_32x32_tb; 

architecture tb of registro_32x32_tb is
    signal 
begin

end tb ; -- tb